module AC_RECEIVER

endmodule