module AC_RECEIVER(
		input			clk
	)

endmodule